
module test(

    );
    reg clk;
    reg reset;
    wire [31:0] WriteData, DataAdr;
    wire MemWrite;

 // instantiate device to be tested
 top_tb dut(clk, reset, WriteData, DataAdr, MemWrite);
 
 // initialize test
 initial
     begin
     reset <= 1; # 22; reset <= 0;
     end
 
 // generate clock to sequence tests
 always
     begin
     clk <= 1; # 5; clk <= 0; # 5;
     end
 
 always @(negedge clk)
 begin
//    $display(" RISCV Simulation Begins!!!!!!");
     if(MemWrite) begin
         if(DataAdr === 7 & WriteData === 32'h05ff_05ff) begin
             $display("Simulation succeeded");
             $stop;
         end 
//         else if (DataAdr !== 34) begin
//             $display("Simulation failed");
//             $stop;
//         end
     end
//     $display(" RISCV Simulation ENDS!!!!!!");
 end
 
////  check results
// always @(negedge clk)
// begin
//    $display(" RISCV Simulation Begins!!!!!!");
//     if(MemWrite) begin
//         if(DataAdr === 100 & WriteData === 25) begin
//             $display("Simulation succeeded");
//             $stop;
//         end 
//         else if (DataAdr !== 96) begin
//             $display("Simulation failed");
//             $stop;
//         end
//     end
//     $display(" RISCV Simulation ENDS!!!!!!");
// end
endmodule
